module ReadyControl(
		input 										st_sts,
		input	 									  mt_wait,
		input 										 mt_ce,
		input 										 st_ce,
		output 										 ready
    );

	always @ (*) begin
		if(st_ce) begin
			if(st_sts)
		
		end
		
	end
	
endmodule
