module dummyRAM(
		input 			 clk,
		input [15: 0]  data,
		input [ 4: 0]  addr,
		
		
    );


endmodule
