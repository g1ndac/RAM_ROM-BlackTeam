module RAM_Controller_Automaton RAM_Controller_Automaton(
		input 													clk,
		input 													rst,
		input 											inAddress,
		inout 												inData,
		input 										  outAddress,
		inout 											  outData,
		output 										  chipEnable,
		output 										outputEnable,
		output 										 writeEnable
		);
		
		

endmodule
